module RISCV_TOP (
	//General Signals
	input wire CLK,
	input wire RSTn,

	//I-Memory Signals
	output wire I_MEM_CSN,
	input wire [31:0] I_MEM_DI,//input from IM
	output reg [11:0] I_MEM_ADDR,//in byte address

	//D-Memory Signals
	output wire D_MEM_CSN,
	input wire [31:0] D_MEM_DI,
	output wire [31:0] D_MEM_DOUT,
	output wire [11:0] D_MEM_ADDR,//in word address
	output wire D_MEM_WEN,
	output wire [3:0] D_MEM_BE,

	//RegFile Signals
	output wire RF_WE,
	output wire [4:0] RF_RA1,
	output wire [4:0] RF_RA2,
	output wire [4:0] RF_WA1,
	input wire [31:0] RF_RD1,
	input wire [31:0] RF_RD2,
	output wire [31:0] RF_WD,
	output wire HALT,                   // if set, terminate program
	output reg [31:0] NUM_INST,         // number of instruction completed
	output wire [31:0] OUTPUT_PORT      // equal RF_WD this port is used for test
	);

	assign OUTPUT_PORT = RF_WD;


/*
	// New added from me
	reg [31:0] PC;
	wire [31:0] NXT_PC;

	assign NXT_PC = (~RSTn) ? 0 :
					(~TAKEN) ? PC + 4 :
					(JUMP_SRC) ? TODO : TODO;

	always @(posedge CLK) begin
		PC <= NXT_PC;
	end
*/


	initial begin
		NUM_INST <= 0;
	end

	// Only allow for NUM_INST
	always @ (negedge CLK) begin
		if (RSTn) begin
			I_MEM_CSN = 0;
			D_MEM_CSN = 0;
		end
		else begin
			I_MEM_CSN = 1;
			D_MEM_CSN = 1;
		end
		if (RSTn) NUM_INST <= NUM_INST + 1;
	end

	// TODO: implement

endmodule //
